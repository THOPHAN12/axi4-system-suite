library verilog;
use verilog.vl_types.all;
entity AXI_Interconnect_Full is
    generic(
        Masters_Num     : integer := 2;
        Slaves_ID_Size  : vl_notype;
        Address_width   : integer := 32;
        S00_Aw_len      : integer := 8;
        S00_Write_data_bus_width: integer := 32;
        S00_Write_data_bytes_num: vl_notype;
        S00_AR_len      : integer := 8;
        S00_Read_data_bus_width: integer := 32;
        S01_Aw_len      : integer := 8;
        S01_AR_len      : integer := 8;
        S01_Write_data_bus_width: integer := 32;
        AXI4_Aw_len     : integer := 8;
        M00_Aw_len      : integer := 8;
        M00_Write_data_bus_width: integer := 32;
        M00_Write_data_bytes_num: vl_notype;
        M00_AR_len      : integer := 8;
        M00_Read_data_bus_width: integer := 32;
        M01_Aw_len      : integer := 8;
        M01_AR_len      : integer := 8;
        M02_Aw_len      : integer := 8;
        M02_AR_len      : integer := 8;
        M02_Read_data_bus_width: integer := 32;
        M03_Aw_len      : integer := 8;
        M03_AR_len      : integer := 8;
        M03_Read_data_bus_width: integer := 32;
        Is_Master_AXI_4 : integer := 1;
        M1_ID           : integer := 0;
        M2_ID           : integer := 1;
        Resp_ID_width   : integer := 2;
        Num_Of_Masters  : integer := 2;
        Num_Of_Slaves   : integer := 4;
        Master_ID_Width : vl_notype;
        AXI4_AR_len     : integer := 8
    );
    port(
        S01_ACLK        : in     vl_logic;
        S01_ARESETN     : in     vl_logic;
        S01_AXI_awaddr  : in     vl_logic_vector;
        S01_AXI_awlen   : in     vl_logic_vector;
        S01_AXI_awsize  : in     vl_logic_vector(2 downto 0);
        S01_AXI_awburst : in     vl_logic_vector(1 downto 0);
        S01_AXI_awlock  : in     vl_logic_vector(1 downto 0);
        S01_AXI_awcache : in     vl_logic_vector(3 downto 0);
        S01_AXI_awprot  : in     vl_logic_vector(2 downto 0);
        S01_AXI_awqos   : in     vl_logic_vector(3 downto 0);
        S01_AXI_awvalid : in     vl_logic;
        S01_AXI_awready : out    vl_logic;
        S01_AXI_wdata   : in     vl_logic_vector;
        S01_AXI_wstrb   : in     vl_logic_vector;
        S01_AXI_wlast   : in     vl_logic;
        S01_AXI_wvalid  : in     vl_logic;
        S01_AXI_wready  : out    vl_logic;
        S01_AXI_bresp   : out    vl_logic_vector(1 downto 0);
        S01_AXI_bvalid  : out    vl_logic;
        S01_AXI_bready  : in     vl_logic;
        S01_AXI_araddr  : in     vl_logic_vector;
        S01_AXI_arlen   : in     vl_logic_vector;
        S01_AXI_arsize  : in     vl_logic_vector(2 downto 0);
        S01_AXI_arburst : in     vl_logic_vector(1 downto 0);
        S01_AXI_arlock  : in     vl_logic_vector(1 downto 0);
        S01_AXI_arcache : in     vl_logic_vector(3 downto 0);
        S01_AXI_arprot  : in     vl_logic_vector(2 downto 0);
        S01_AXI_arregion: in     vl_logic_vector(3 downto 0);
        S01_AXI_arqos   : in     vl_logic_vector(3 downto 0);
        S01_AXI_arvalid : in     vl_logic;
        S01_AXI_arready : out    vl_logic;
        S01_AXI_rdata   : out    vl_logic_vector;
        S01_AXI_rresp   : out    vl_logic_vector(1 downto 0);
        S01_AXI_rlast   : out    vl_logic;
        S01_AXI_rvalid  : out    vl_logic;
        S01_AXI_rready  : in     vl_logic;
        ACLK            : in     vl_logic;
        ARESETN         : in     vl_logic;
        S00_ACLK        : in     vl_logic;
        S00_ARESETN     : in     vl_logic;
        S00_AXI_awaddr  : in     vl_logic_vector;
        S00_AXI_awlen   : in     vl_logic_vector;
        S00_AXI_awsize  : in     vl_logic_vector(2 downto 0);
        S00_AXI_awburst : in     vl_logic_vector(1 downto 0);
        S00_AXI_awlock  : in     vl_logic_vector(1 downto 0);
        S00_AXI_awcache : in     vl_logic_vector(3 downto 0);
        S00_AXI_awprot  : in     vl_logic_vector(2 downto 0);
        S00_AXI_awqos   : in     vl_logic_vector(3 downto 0);
        S00_AXI_awvalid : in     vl_logic;
        S00_AXI_awready : out    vl_logic;
        S00_AXI_wdata   : in     vl_logic_vector;
        S00_AXI_wstrb   : in     vl_logic_vector;
        S00_AXI_wlast   : in     vl_logic;
        S00_AXI_wvalid  : in     vl_logic;
        S00_AXI_wready  : out    vl_logic;
        S00_AXI_bresp   : out    vl_logic_vector(1 downto 0);
        S00_AXI_bvalid  : out    vl_logic;
        S00_AXI_bready  : in     vl_logic;
        S00_AXI_araddr  : in     vl_logic_vector;
        S00_AXI_arlen   : in     vl_logic_vector;
        S00_AXI_arsize  : in     vl_logic_vector(2 downto 0);
        S00_AXI_arburst : in     vl_logic_vector(1 downto 0);
        S00_AXI_arlock  : in     vl_logic_vector(1 downto 0);
        S00_AXI_arcache : in     vl_logic_vector(3 downto 0);
        S00_AXI_arprot  : in     vl_logic_vector(2 downto 0);
        S00_AXI_arregion: in     vl_logic_vector(3 downto 0);
        S00_AXI_arqos   : in     vl_logic_vector(3 downto 0);
        S00_AXI_arvalid : in     vl_logic;
        S00_AXI_arready : out    vl_logic;
        S00_AXI_rdata   : out    vl_logic_vector;
        S00_AXI_rresp   : out    vl_logic_vector(1 downto 0);
        S00_AXI_rlast   : out    vl_logic;
        S00_AXI_rvalid  : out    vl_logic;
        S00_AXI_rready  : in     vl_logic;
        M00_ACLK        : in     vl_logic;
        M00_ARESETN     : in     vl_logic;
        M00_AXI_awaddr_ID: out    vl_logic_vector;
        M00_AXI_awaddr  : out    vl_logic_vector;
        M00_AXI_awlen   : out    vl_logic_vector;
        M00_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M00_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M00_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M00_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M00_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M00_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M00_AXI_awvalid : out    vl_logic;
        M00_AXI_awready : in     vl_logic;
        M00_AXI_wdata   : out    vl_logic_vector;
        M00_AXI_wstrb   : out    vl_logic_vector;
        M00_AXI_wlast   : out    vl_logic;
        M00_AXI_wvalid  : out    vl_logic;
        M00_AXI_wready  : in     vl_logic;
        M00_AXI_BID     : in     vl_logic_vector;
        M00_AXI_bresp   : in     vl_logic_vector(1 downto 0);
        M00_AXI_bvalid  : in     vl_logic;
        M00_AXI_bready  : out    vl_logic;
        M00_AXI_araddr  : out    vl_logic_vector;
        M00_AXI_arlen   : out    vl_logic_vector;
        M00_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M00_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M00_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M00_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M00_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M00_AXI_arvalid : out    vl_logic;
        M00_AXI_arready : in     vl_logic;
        M00_AXI_rdata   : in     vl_logic_vector;
        M00_AXI_rresp   : in     vl_logic_vector(1 downto 0);
        M00_AXI_rlast   : in     vl_logic;
        M00_AXI_rvalid  : in     vl_logic;
        M00_AXI_rready  : out    vl_logic;
        M01_ACLK        : in     vl_logic;
        M01_ARESETN     : in     vl_logic;
        M01_AXI_awaddr_ID: out    vl_logic_vector;
        M01_AXI_awaddr  : out    vl_logic_vector;
        M01_AXI_awlen   : out    vl_logic_vector;
        M01_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_awvalid : out    vl_logic;
        M01_AXI_awready : in     vl_logic;
        M01_AXI_wdata   : out    vl_logic_vector;
        M01_AXI_wstrb   : out    vl_logic_vector;
        M01_AXI_wlast   : out    vl_logic;
        M01_AXI_wvalid  : out    vl_logic;
        M01_AXI_wready  : in     vl_logic;
        M01_AXI_BID     : in     vl_logic_vector;
        M01_AXI_bresp   : in     vl_logic_vector(1 downto 0);
        M01_AXI_bvalid  : in     vl_logic;
        M01_AXI_bready  : out    vl_logic;
        M01_AXI_araddr  : out    vl_logic_vector;
        M01_AXI_arlen   : out    vl_logic_vector;
        M01_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M01_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_arvalid : out    vl_logic;
        M01_AXI_arready : in     vl_logic;
        M01_AXI_rdata   : in     vl_logic_vector;
        M01_AXI_rresp   : in     vl_logic_vector(1 downto 0);
        M01_AXI_rlast   : in     vl_logic;
        M01_AXI_rvalid  : in     vl_logic;
        M01_AXI_rready  : out    vl_logic;
        slave0_addr1    : in     vl_logic_vector(31 downto 0);
        slave0_addr2    : in     vl_logic_vector(31 downto 0);
        slave1_addr1    : in     vl_logic_vector(31 downto 0);
        slave1_addr2    : in     vl_logic_vector(31 downto 0);
        slave2_addr1    : in     vl_logic_vector(31 downto 0);
        slave2_addr2    : in     vl_logic_vector(31 downto 0);
        slave3_addr1    : in     vl_logic_vector(31 downto 0);
        slave3_addr2    : in     vl_logic_vector(31 downto 0);
        M02_ACLK        : in     vl_logic;
        M02_ARESETN     : in     vl_logic;
        M02_AXI_araddr  : out    vl_logic_vector;
        M02_AXI_arlen   : out    vl_logic_vector;
        M02_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M02_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M02_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M02_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M02_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M02_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M02_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M02_AXI_arvalid : out    vl_logic;
        M02_AXI_arready : in     vl_logic;
        M02_AXI_rdata   : in     vl_logic_vector;
        M02_AXI_rresp   : in     vl_logic_vector(1 downto 0);
        M02_AXI_rlast   : in     vl_logic;
        M02_AXI_rvalid  : in     vl_logic;
        M02_AXI_rready  : out    vl_logic;
        M03_ACLK        : in     vl_logic;
        M03_ARESETN     : in     vl_logic;
        M03_AXI_araddr  : out    vl_logic_vector;
        M03_AXI_arlen   : out    vl_logic_vector;
        M03_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M03_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M03_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M03_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M03_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M03_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M03_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M03_AXI_arvalid : out    vl_logic;
        M03_AXI_arready : in     vl_logic;
        M03_AXI_rdata   : in     vl_logic_vector;
        M03_AXI_rresp   : in     vl_logic_vector(1 downto 0);
        M03_AXI_rlast   : in     vl_logic;
        M03_AXI_rvalid  : in     vl_logic;
        M03_AXI_rready  : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of Masters_Num : constant is 1;
    attribute mti_svvh_generic_type of Slaves_ID_Size : constant is 3;
    attribute mti_svvh_generic_type of Address_width : constant is 1;
    attribute mti_svvh_generic_type of S00_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of S00_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of S00_Write_data_bytes_num : constant is 3;
    attribute mti_svvh_generic_type of S00_AR_len : constant is 1;
    attribute mti_svvh_generic_type of S00_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of S01_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of S01_AR_len : constant is 1;
    attribute mti_svvh_generic_type of S01_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of AXI4_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of M00_Write_data_bytes_num : constant is 3;
    attribute mti_svvh_generic_type of M00_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of M01_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M01_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M02_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M02_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M02_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of M03_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M03_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M03_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of Is_Master_AXI_4 : constant is 1;
    attribute mti_svvh_generic_type of M1_ID : constant is 1;
    attribute mti_svvh_generic_type of M2_ID : constant is 1;
    attribute mti_svvh_generic_type of Resp_ID_width : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Masters : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Slaves : constant is 1;
    attribute mti_svvh_generic_type of Master_ID_Width : constant is 3;
    attribute mti_svvh_generic_type of AXI4_AR_len : constant is 1;
end AXI_Interconnect_Full;
