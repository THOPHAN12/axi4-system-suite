library verilog;
use verilog.vl_types.all;
entity test_case2 is
end test_case2;
