library verilog;
use verilog.vl_types.all;
entity test_case4 is
end test_case4;
