library verilog;
use verilog.vl_types.all;
entity alu_master_system is
    generic(
        ADDR_WIDTH      : integer := 32;
        DATA_WIDTH      : integer := 32;
        ID_WIDTH        : integer := 4;
        MEM_SIZE        : integer := 256;
        Masters_Num     : integer := 2;
        Slaves_ID_Size  : integer := 1;
        Address_width   : integer := 32;
        S00_Aw_len      : integer := 8;
        S00_Write_data_bus_width: integer := 32;
        S00_Write_data_bytes_num: integer := 4;
        S00_AR_len      : integer := 8;
        S00_Read_data_bus_width: integer := 32;
        S01_Aw_len      : integer := 8;
        S01_Write_data_bus_width: integer := 32;
        S01_AR_len      : integer := 8;
        M00_Aw_len      : integer := 8;
        M00_Write_data_bus_width: integer := 32;
        M00_Write_data_bytes_num: integer := 4;
        M00_AR_len      : integer := 8;
        M00_Read_data_bus_width: integer := 32;
        M01_Aw_len      : integer := 8;
        M01_AR_len      : integer := 8;
        M02_Aw_len      : integer := 8;
        M02_AR_len      : integer := 8;
        M02_Read_data_bus_width: integer := 32;
        M03_Aw_len      : integer := 8;
        M03_AR_len      : integer := 8;
        M03_Read_data_bus_width: integer := 32;
        Is_Master_AXI_4 : vl_logic := Hi1;
        M1_ID           : integer := 0;
        M2_ID           : integer := 1;
        Resp_ID_width   : integer := 2;
        Num_Of_Masters  : integer := 2;
        Num_Of_Slaves   : integer := 4;
        Master_ID_Width : integer := 1;
        AXI4_AR_len     : integer := 8;
        AXI4_Aw_len     : integer := 8;
        SLAVE0_ADDR1    : integer := 0;
        SLAVE0_ADDR2    : integer := 1073741823;
        SLAVE1_ADDR1    : integer := 1073741824;
        SLAVE1_ADDR2    : integer := 2147483647;
        SLAVE2_ADDR1    : vl_logic_vector(31 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SLAVE2_ADDR2    : vl_logic_vector(31 downto 0) := (Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        SLAVE3_ADDR1    : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SLAVE3_ADDR2    : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1)
    );
    port(
        ACLK            : in     vl_logic;
        ARESETN         : in     vl_logic;
        master0_start   : in     vl_logic;
        master0_busy    : out    vl_logic;
        master0_done    : out    vl_logic;
        master1_start   : in     vl_logic;
        master1_busy    : out    vl_logic;
        master1_done    : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_SIZE : constant is 1;
    attribute mti_svvh_generic_type of Masters_Num : constant is 1;
    attribute mti_svvh_generic_type of Slaves_ID_Size : constant is 1;
    attribute mti_svvh_generic_type of Address_width : constant is 1;
    attribute mti_svvh_generic_type of S00_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of S00_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of S00_Write_data_bytes_num : constant is 1;
    attribute mti_svvh_generic_type of S00_AR_len : constant is 1;
    attribute mti_svvh_generic_type of S00_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of S01_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of S01_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of S01_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Write_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of M00_Write_data_bytes_num : constant is 1;
    attribute mti_svvh_generic_type of M00_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of M01_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M01_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M02_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M02_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M02_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of M03_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M03_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M03_Read_data_bus_width : constant is 1;
    attribute mti_svvh_generic_type of Is_Master_AXI_4 : constant is 1;
    attribute mti_svvh_generic_type of M1_ID : constant is 1;
    attribute mti_svvh_generic_type of M2_ID : constant is 1;
    attribute mti_svvh_generic_type of Resp_ID_width : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Masters : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Slaves : constant is 1;
    attribute mti_svvh_generic_type of Master_ID_Width : constant is 1;
    attribute mti_svvh_generic_type of AXI4_AR_len : constant is 1;
    attribute mti_svvh_generic_type of AXI4_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of SLAVE0_ADDR1 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE0_ADDR2 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE1_ADDR1 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE1_ADDR2 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE2_ADDR1 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE2_ADDR2 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE3_ADDR1 : constant is 1;
    attribute mti_svvh_generic_type of SLAVE3_ADDR2 : constant is 1;
end alu_master_system;
