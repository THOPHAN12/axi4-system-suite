library verilog;
use verilog.vl_types.all;
entity Write_Addr_Channel_Dec is
    generic(
        Num_OF_Masters  : integer := 2;
        Masters_ID_Size : vl_notype;
        Address_width   : integer := 32;
        AXI4_Aw_len     : integer := 8;
        Num_Of_Slaves   : integer := 4;
        Base_Addr_Width : vl_notype
    );
    port(
        Master_AXI_awaddr_ID: in     vl_logic_vector;
        Master_AXI_awaddr: in     vl_logic_vector;
        Master_AXI_awlen: in     vl_logic_vector;
        Master_AXI_awsize: in     vl_logic_vector(2 downto 0);
        Master_AXI_awburst: in     vl_logic_vector(1 downto 0);
        Master_AXI_awlock: in     vl_logic_vector(1 downto 0);
        Master_AXI_awcache: in     vl_logic_vector(3 downto 0);
        Master_AXI_awprot: in     vl_logic_vector(2 downto 0);
        Master_AXI_awqos: in     vl_logic_vector(3 downto 0);
        Master_AXI_awvalid: in     vl_logic;
        M00_AXI_awaddr_ID: out    vl_logic_vector;
        M00_AXI_awaddr  : out    vl_logic_vector;
        M00_AXI_awlen   : out    vl_logic_vector;
        M00_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M00_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M00_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M00_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M00_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M00_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M00_AXI_awvalid : out    vl_logic;
        M00_AXI_awready : in     vl_logic;
        M01_AXI_awaddr_ID: out    vl_logic_vector;
        M01_AXI_awaddr  : out    vl_logic_vector;
        M01_AXI_awlen   : out    vl_logic_vector;
        M01_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_awvalid : out    vl_logic;
        M01_AXI_awready : in     vl_logic;
        M02_AXI_awaddr_ID: out    vl_logic_vector;
        M02_AXI_awaddr  : out    vl_logic_vector;
        M02_AXI_awlen   : out    vl_logic_vector;
        M02_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M02_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M02_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M02_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M02_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M02_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M02_AXI_awvalid : out    vl_logic;
        M02_AXI_awready : in     vl_logic;
        M03_AXI_awaddr_ID: out    vl_logic_vector;
        M03_AXI_awaddr  : out    vl_logic_vector;
        M03_AXI_awlen   : out    vl_logic_vector;
        M03_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M03_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M03_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M03_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M03_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M03_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M03_AXI_awvalid : out    vl_logic;
        M03_AXI_awready : in     vl_logic;
        Sel_Slave_Ready : out    vl_logic;
        Q_Enables       : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of Num_OF_Masters : constant is 1;
    attribute mti_svvh_generic_type of Masters_ID_Size : constant is 3;
    attribute mti_svvh_generic_type of Address_width : constant is 1;
    attribute mti_svvh_generic_type of AXI4_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Slaves : constant is 1;
    attribute mti_svvh_generic_type of Base_Addr_Width : constant is 3;
end Write_Addr_Channel_Dec;
