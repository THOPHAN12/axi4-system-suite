library verilog;
use verilog.vl_types.all;
entity test_case1_read is
end test_case1_read;
