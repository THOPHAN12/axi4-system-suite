library verilog;
use verilog.vl_types.all;
entity AXI_Interconnect is
    port(
        G_clk           : in     vl_logic;
        G_reset         : in     vl_logic;
        M0_RREADY       : in     vl_logic;
        M0_ARADDR       : in     vl_logic_vector(31 downto 0);
        M0_ARLEN        : in     vl_logic_vector(3 downto 0);
        M0_ARSIZE       : in     vl_logic_vector(2 downto 0);
        M0_ARBURST      : in     vl_logic_vector(1 downto 0);
        M0_ARVALID      : in     vl_logic;
        M1_RREADY       : in     vl_logic;
        M1_ARADDR       : in     vl_logic_vector(31 downto 0);
        M1_ARLEN        : in     vl_logic_vector(3 downto 0);
        M1_ARSIZE       : in     vl_logic_vector(2 downto 0);
        M1_ARBURST      : in     vl_logic_vector(1 downto 0);
        M1_ARVALID      : in     vl_logic;
        S0_ARREADY      : in     vl_logic;
        S0_RVALID       : in     vl_logic;
        S0_RLAST        : in     vl_logic;
        S0_RRESP        : in     vl_logic_vector(1 downto 0);
        S0_RDATA        : in     vl_logic_vector(31 downto 0);
        S1_ARREADY      : in     vl_logic;
        S1_RVALID       : in     vl_logic;
        S1_RLAST        : in     vl_logic;
        S1_RRESP        : in     vl_logic_vector(1 downto 0);
        S1_RDATA        : in     vl_logic_vector(31 downto 0);
        slave0_addr1    : in     vl_logic_vector(31 downto 0);
        slave0_addr2    : in     vl_logic_vector(31 downto 0);
        slave1_addr1    : in     vl_logic_vector(31 downto 0);
        slave1_addr2    : in     vl_logic_vector(31 downto 0);
        ARREADY_M0      : out    vl_logic;
        RVALID_M0       : out    vl_logic;
        RLAST_M0        : out    vl_logic;
        RRESP_M0        : out    vl_logic_vector(1 downto 0);
        RDATA_M0        : out    vl_logic_vector(31 downto 0);
        ARREADY_M1      : out    vl_logic;
        RVALID_M1       : out    vl_logic;
        RLAST_M1        : out    vl_logic;
        RRESP_M1        : out    vl_logic_vector(1 downto 0);
        RDATA_M1        : out    vl_logic_vector(31 downto 0);
        ARADDR_S0       : out    vl_logic_vector(31 downto 0);
        ARLEN_S0        : out    vl_logic_vector(3 downto 0);
        ARSIZE_S0       : out    vl_logic_vector(2 downto 0);
        ARBURST_S0      : out    vl_logic_vector(1 downto 0);
        ARVALID_S0      : out    vl_logic;
        RREADY_S0       : out    vl_logic;
        ARADDR_S1       : out    vl_logic_vector(31 downto 0);
        ARLEN_S1        : out    vl_logic_vector(3 downto 0);
        ARSIZE_S1       : out    vl_logic_vector(2 downto 0);
        ARBURST_S1      : out    vl_logic_vector(1 downto 0);
        ARVALID_S1      : out    vl_logic;
        RREADY_S1       : out    vl_logic
    );
end AXI_Interconnect;
