library verilog;
use verilog.vl_types.all;
entity test_case3 is
end test_case3;
