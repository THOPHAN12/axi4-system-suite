library verilog;
use verilog.vl_types.all;
entity AR_Channel_Controller_Top is
    generic(
        Masters_Num     : integer := 2;
        Slaves_ID_Size  : vl_notype;
        Address_width   : integer := 32;
        S00_AR_len      : integer := 8;
        S01_AR_len      : integer := 8;
        M00_AR_len      : integer := 8;
        M01_AR_len      : integer := 8;
        M02_AR_len      : integer := 8;
        M03_AR_len      : integer := 8;
        AXI4_AR_len     : integer := 8;
        Num_Of_Slaves   : integer := 4
    );
    port(
        AR_Access_Grant : out    vl_logic;
        AR_Selected_Slave: out    vl_logic_vector;
        AR_Channel_Request: out    vl_logic;
        ACLK            : in     vl_logic;
        ARESETN         : in     vl_logic;
        S00_ACLK        : in     vl_logic;
        S00_ARESETN     : in     vl_logic;
        S00_AXI_araddr  : in     vl_logic_vector;
        S00_AXI_arlen   : in     vl_logic_vector;
        S00_AXI_arsize  : in     vl_logic_vector(2 downto 0);
        S00_AXI_arburst : in     vl_logic_vector(1 downto 0);
        S00_AXI_arlock  : in     vl_logic_vector(1 downto 0);
        S00_AXI_arcache : in     vl_logic_vector(3 downto 0);
        S00_AXI_arprot  : in     vl_logic_vector(2 downto 0);
        S00_AXI_arqos   : in     vl_logic_vector(3 downto 0);
        S00_AXI_arregion: in     vl_logic_vector(3 downto 0);
        S00_AXI_arvalid : in     vl_logic;
        S00_AXI_arready : out    vl_logic;
        S01_ACLK        : in     vl_logic;
        S01_ARESETN     : in     vl_logic;
        S01_AXI_araddr  : in     vl_logic_vector;
        S01_AXI_arlen   : in     vl_logic_vector;
        S01_AXI_arsize  : in     vl_logic_vector(2 downto 0);
        S01_AXI_arburst : in     vl_logic_vector(1 downto 0);
        S01_AXI_arlock  : in     vl_logic_vector(1 downto 0);
        S01_AXI_arcache : in     vl_logic_vector(3 downto 0);
        S01_AXI_arprot  : in     vl_logic_vector(2 downto 0);
        S01_AXI_arqos   : in     vl_logic_vector(3 downto 0);
        S01_AXI_arregion: in     vl_logic_vector(3 downto 0);
        S01_AXI_arvalid : in     vl_logic;
        S01_AXI_arready : out    vl_logic;
        M00_ACLK        : in     vl_logic;
        M00_ARESETN     : in     vl_logic;
        M00_AXI_araddr_ID: out    vl_logic_vector;
        M00_AXI_araddr  : out    vl_logic_vector;
        M00_AXI_arlen   : out    vl_logic_vector;
        M00_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M00_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M00_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M00_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M00_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M00_AXI_arvalid : out    vl_logic;
        M00_AXI_arready : in     vl_logic;
        M01_ACLK        : in     vl_logic;
        M01_ARESETN     : in     vl_logic;
        M01_AXI_araddr_ID: out    vl_logic_vector;
        M01_AXI_araddr  : out    vl_logic_vector;
        M01_AXI_arlen   : out    vl_logic_vector;
        M01_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M01_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_arvalid : out    vl_logic;
        M01_AXI_arready : in     vl_logic;
        M02_ACLK        : in     vl_logic;
        M02_ARESETN     : in     vl_logic;
        M02_AXI_araddr_ID: out    vl_logic_vector;
        M02_AXI_araddr  : out    vl_logic_vector;
        M02_AXI_arlen   : out    vl_logic_vector;
        M02_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M02_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M02_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M02_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M02_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M02_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M02_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M02_AXI_arvalid : out    vl_logic;
        M02_AXI_arready : in     vl_logic;
        M03_ACLK        : in     vl_logic;
        M03_ARESETN     : in     vl_logic;
        M03_AXI_araddr_ID: out    vl_logic_vector;
        M03_AXI_araddr  : out    vl_logic_vector;
        M03_AXI_arlen   : out    vl_logic_vector;
        M03_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M03_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M03_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M03_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M03_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M03_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M03_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M03_AXI_arvalid : out    vl_logic;
        M03_AXI_arready : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of Masters_Num : constant is 1;
    attribute mti_svvh_generic_type of Slaves_ID_Size : constant is 3;
    attribute mti_svvh_generic_type of Address_width : constant is 1;
    attribute mti_svvh_generic_type of S00_AR_len : constant is 1;
    attribute mti_svvh_generic_type of S01_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M00_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M01_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M02_AR_len : constant is 1;
    attribute mti_svvh_generic_type of M03_AR_len : constant is 1;
    attribute mti_svvh_generic_type of AXI4_AR_len : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Slaves : constant is 1;
end AR_Channel_Controller_Top;
