library verilog;
use verilog.vl_types.all;
entity BReady_MUX_2_1_tb is
end BReady_MUX_2_1_tb;
