library verilog;
use verilog.vl_types.all;
entity test_case1 is
end test_case1;
