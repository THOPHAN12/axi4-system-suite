`timescale 1ns/1ps

interface bready_mux_if ();
    logic select;
    logic m0_ready;
    logic m1_ready;
    logic sel_ready;
endinterface

