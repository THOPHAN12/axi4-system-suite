library verilog;
use verilog.vl_types.all;
entity AW_Channel_Controller_Top is
    generic(
        Masters_Num     : integer := 2;
        Slaves_ID_Size  : vl_notype;
        Address_width   : integer := 32;
        S00_Aw_len      : integer := 8;
        S01_Aw_len      : integer := 8;
        Is_Master_AXI_4 : integer := 1;
        AXI4_Aw_len     : integer := 8;
        M00_Aw_len      : integer := 8;
        M01_Aw_len      : integer := 8;
        Num_Of_Slaves   : integer := 2
    );
    port(
        AW_Access_Grant : out    vl_logic;
        AW_Selected_Slave: out    vl_logic_vector;
        Queue_Is_Full   : in     vl_logic;
        Token           : out    vl_logic;
        \Rem\           : out    vl_logic_vector;
        Num_Of_Compl_Bursts: out    vl_logic_vector;
        Load_The_Original_Signals: out    vl_logic;
        ACLK            : in     vl_logic;
        ARESETN         : in     vl_logic;
        S00_ACLK        : in     vl_logic;
        S00_ARESETN     : in     vl_logic;
        S00_AXI_awaddr  : in     vl_logic_vector;
        S00_AXI_awlen   : in     vl_logic_vector;
        S00_AXI_awsize  : in     vl_logic_vector(2 downto 0);
        S00_AXI_awburst : in     vl_logic_vector(1 downto 0);
        S00_AXI_awlock  : in     vl_logic_vector(1 downto 0);
        S00_AXI_awcache : in     vl_logic_vector(3 downto 0);
        S00_AXI_awprot  : in     vl_logic_vector(2 downto 0);
        S00_AXI_awqos   : in     vl_logic_vector(3 downto 0);
        S00_AXI_awvalid : in     vl_logic;
        S00_AXI_awready : out    vl_logic;
        S01_ACLK        : in     vl_logic;
        S01_ARESETN     : in     vl_logic;
        S01_AXI_awaddr  : in     vl_logic_vector;
        S01_AXI_awlen   : in     vl_logic_vector;
        S01_AXI_awsize  : in     vl_logic_vector(2 downto 0);
        S01_AXI_awburst : in     vl_logic_vector(1 downto 0);
        S01_AXI_awlock  : in     vl_logic_vector(1 downto 0);
        S01_AXI_awcache : in     vl_logic_vector(3 downto 0);
        S01_AXI_awprot  : in     vl_logic_vector(2 downto 0);
        S01_AXI_awqos   : in     vl_logic_vector(3 downto 0);
        S01_AXI_awvalid : in     vl_logic;
        S01_AXI_awready : out    vl_logic;
        M00_ACLK        : in     vl_logic;
        M00_ARESETN     : in     vl_logic;
        M00_AXI_awaddr_ID: out    vl_logic_vector;
        M00_AXI_awaddr  : out    vl_logic_vector;
        M00_AXI_awlen   : out    vl_logic_vector;
        M00_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M00_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M00_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M00_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M00_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M00_AXI_awvalid : out    vl_logic;
        M00_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M00_AXI_awready : in     vl_logic;
        M01_ACLK        : in     vl_logic;
        M01_ARESETN     : in     vl_logic;
        M01_AXI_awaddr_ID: out    vl_logic_vector;
        M01_AXI_awaddr  : out    vl_logic_vector;
        M01_AXI_awlen   : out    vl_logic_vector;
        M01_AXI_awsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_awburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_awlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_awcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_awprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_awvalid : out    vl_logic;
        M01_AXI_awqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_awready : in     vl_logic;
        Q_Enable_W_Data : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of Masters_Num : constant is 1;
    attribute mti_svvh_generic_type of Slaves_ID_Size : constant is 3;
    attribute mti_svvh_generic_type of Address_width : constant is 1;
    attribute mti_svvh_generic_type of S00_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of S01_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of Is_Master_AXI_4 : constant is 1;
    attribute mti_svvh_generic_type of AXI4_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M00_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of M01_Aw_len : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Slaves : constant is 1;
end AW_Channel_Controller_Top;
