library verilog;
use verilog.vl_types.all;
entity test_case5 is
end test_case5;
