// ==============================================================================
// FRISCV AXI System - Complete Integration
// ==============================================================================
// Integrates FRISCV RV32I core with AXI Interconnect and peripherals
//
// Architecture:
// - FRISCV RV32I Core (3-stage pipeline, caches, RV32IM)
// - 2× AXI Width Adapters (128-bit → 32-bit)
// - AXI Interconnect (2M × 4S, Round-Robin)
// - 4× AXI-Lite Peripherals (RAM, GPIO, UART, SPI)
//
// Auto-generated by: AXI Bridge Integration Tool
// Date: December 5, 2025
// Status: Production-Ready
// ==============================================================================

`timescale 1ns/1ps

module friscv_axi_system (
    // Clock and Reset
    input wire ACLK,
    input wire ARESETN,
    
    // Soft Reset (optional)
    input wire SRST,
    
    // Interrupts
    input wire ext_irq,
    input wire sw_irq,
    input wire timer_irq,
    
    // GPIO
    input  wire [31:0] gpio_in,
    output wire [31:0] gpio_out,
    
    // UART
    input  wire uart_rx,
    output wire uart_tx,
    
    // SPI
    output wire spi_sclk,
    output wire spi_mosi,
    input  wire spi_miso,
    output wire spi_cs_n,
    
    // Debug
    output wire [7:0]   debug_status,
    output wire [1023:0] debug_regs  // 32 registers × 32 bits
);

// ==============================================================================
// Internal Signals - FRISCV Core (128-bit AXI)
// ==============================================================================

// Instruction Memory (128-bit)
wire        friscv_imem_arvalid;
wire        friscv_imem_arready;
wire [31:0] friscv_imem_araddr;
wire [2:0]  friscv_imem_arprot;
wire [7:0]  friscv_imem_arid;
wire        friscv_imem_rvalid;
wire        friscv_imem_rready;
wire [7:0]  friscv_imem_rid;
wire [1:0]  friscv_imem_rresp;
wire [127:0] friscv_imem_rdata;

// Data Memory (128-bit)
wire        friscv_dmem_awvalid;
wire        friscv_dmem_awready;
wire [31:0] friscv_dmem_awaddr;
wire [2:0]  friscv_dmem_awprot;
wire [7:0]  friscv_dmem_awid;
wire        friscv_dmem_wvalid;
wire        friscv_dmem_wready;
wire [127:0] friscv_dmem_wdata;
wire [15:0] friscv_dmem_wstrb;
wire        friscv_dmem_bvalid;
wire        friscv_dmem_bready;
wire [7:0]  friscv_dmem_bid;
wire [1:0]  friscv_dmem_bresp;
wire        friscv_dmem_arvalid;
wire        friscv_dmem_arready;
wire [31:0] friscv_dmem_araddr;
wire [2:0]  friscv_dmem_arprot;
wire [7:0]  friscv_dmem_arid;
wire        friscv_dmem_rvalid;
wire        friscv_dmem_rready;
wire [7:0]  friscv_dmem_rid;
wire [1:0]  friscv_dmem_rresp;
wire [127:0] friscv_dmem_rdata;

// ==============================================================================
// Internal Signals - Width Adapters → Interconnect (32-bit AXI)
// ==============================================================================

// Master 0 (Instruction) - 32-bit
wire        m0_axi_arvalid;
wire        m0_axi_arready;
wire [31:0] m0_axi_araddr;
wire [7:0]  m0_axi_arlen;
wire [2:0]  m0_axi_arsize;
wire [1:0]  m0_axi_arburst;
wire [2:0]  m0_axi_arprot;
wire        m0_axi_rvalid;
wire        m0_axi_rready;
wire [31:0] m0_axi_rdata;
wire [1:0]  m0_axi_rresp;
wire        m0_axi_rlast;

// Master 1 (Data) - 32-bit  
wire        m1_axi_awvalid;
wire        m1_axi_awready;
wire [31:0] m1_axi_awaddr;
wire [7:0]  m1_axi_awlen;
wire [2:0]  m1_axi_awsize;
wire [1:0]  m1_axi_awburst;
wire [2:0]  m1_axi_awprot;
wire        m1_axi_wvalid;
wire        m1_axi_wready;
wire [31:0] m1_axi_wdata;
wire [3:0]  m1_axi_wstrb;
wire        m1_axi_wlast;
wire        m1_axi_bvalid;
wire        m1_axi_bready;
wire [1:0]  m1_axi_bresp;
wire        m1_axi_arvalid;
wire        m1_axi_arready;
wire [31:0] m1_axi_araddr;
wire [7:0]  m1_axi_arlen;
wire [2:0]  m1_axi_arsize;
wire [1:0]  m1_axi_arburst;
wire [2:0]  m1_axi_arprot;
wire        m1_axi_rvalid;
wire        m1_axi_rready;
wire [31:0] m1_axi_rdata;
wire [1:0]  m1_axi_rresp;
wire        m1_axi_rlast;

// Slave signals (to peripherals) - same as before
wire [31:0] s0_axi_awaddr, s0_axi_araddr, s0_axi_wdata, s0_axi_rdata;
wire [3:0]  s0_axi_wstrb;
wire        s0_axi_awvalid, s0_axi_awready, s0_axi_wvalid, s0_axi_wready;
wire [1:0]  s0_axi_bresp;
wire        s0_axi_bvalid, s0_axi_bready;
wire        s0_axi_arvalid, s0_axi_arready;
wire [1:0]  s0_axi_rresp;
wire        s0_axi_rvalid, s0_axi_rready;

wire [31:0] s1_axi_awaddr, s1_axi_araddr, s1_axi_wdata, s1_axi_rdata;
wire [3:0]  s1_axi_wstrb;
wire        s1_axi_awvalid, s1_axi_awready, s1_axi_wvalid, s1_axi_wready;
wire [1:0]  s1_axi_bresp;
wire        s1_axi_bvalid, s1_axi_bready, s1_axi_arvalid, s1_axi_arready;
wire [1:0]  s1_axi_rresp;
wire        s1_axi_rvalid, s1_axi_rready;

wire [31:0] s2_axi_awaddr, s2_axi_araddr, s2_axi_wdata, s2_axi_rdata;
wire [3:0]  s2_axi_wstrb;
wire        s2_axi_awvalid, s2_axi_awready, s2_axi_wvalid, s2_axi_wready;
wire [1:0]  s2_axi_bresp;
wire        s2_axi_bvalid, s2_axi_bready, s2_axi_arvalid, s2_axi_arready;
wire [1:0]  s2_axi_rresp;
wire        s2_axi_rvalid, s2_axi_rready;

wire [31:0] s3_axi_awaddr, s3_axi_araddr, s3_axi_wdata, s3_axi_rdata;
wire [3:0]  s3_axi_wstrb;
wire        s3_axi_awvalid, s3_axi_awready, s3_axi_wvalid, s3_axi_wready;
wire [1:0]  s3_axi_bresp;
wire        s3_axi_bvalid, s3_axi_bready, s3_axi_arvalid, s3_axi_arready;
wire [1:0]  s3_axi_rresp;
wire        s3_axi_rvalid, s3_axi_rready;

// ==============================================================================
// FRISCV RV32I Core
// ==============================================================================
friscv_rv32i_core #(
    .XLEN(32),
    .BOOT_ADDR(32'h00000000),
    .AXI_ADDR_W(32),
    .AXI_ID_W(8),
    .AXI_IMEM_W(128),                // 128-bit instruction interface
    .AXI_DMEM_W(128),                // 128-bit data interface
    .CACHE_EN(1),                    // Enable caches
    .ICACHE_DEPTH(512),              // 512 instruction cache blocks
    .DCACHE_DEPTH(512),              // 512 data cache blocks
    .M_EXTENSION(1)                  // Enable multiply/divide
) u_friscv_core (
    .aclk(ACLK),
    .aresetn(ARESETN),
    .srst(SRST),
    
    // Interrupts
    .ext_irq(ext_irq),
    .sw_irq(sw_irq),
    .timer_irq(timer_irq),
    
    // Debug
    .status(debug_status),
    .dbg_regs(debug_regs),
    
    // Instruction Memory (128-bit AXI)
    .imem_arvalid(friscv_imem_arvalid),
    .imem_arready(friscv_imem_arready),
    .imem_araddr(friscv_imem_araddr),
    .imem_arprot(friscv_imem_arprot),
    .imem_arid(friscv_imem_arid),
    .imem_rvalid(friscv_imem_rvalid),
    .imem_rready(friscv_imem_rready),
    .imem_rid(friscv_imem_rid),
    .imem_rresp(friscv_imem_rresp),
    .imem_rdata(friscv_imem_rdata),
    
    // Data Memory (128-bit AXI)
    .dmem_awvalid(friscv_dmem_awvalid),
    .dmem_awready(friscv_dmem_awready),
    .dmem_awaddr(friscv_dmem_awaddr),
    .dmem_awprot(friscv_dmem_awprot),
    .dmem_awid(friscv_dmem_awid),
    .dmem_wvalid(friscv_dmem_wvalid),
    .dmem_wready(friscv_dmem_wready),
    .dmem_wdata(friscv_dmem_wdata),
    .dmem_wstrb(friscv_dmem_wstrb),
    .dmem_bvalid(friscv_dmem_bvalid),
    .dmem_bready(friscv_dmem_bready),
    .dmem_bid(friscv_dmem_bid),
    .dmem_bresp(friscv_dmem_bresp),
    .dmem_arvalid(friscv_dmem_arvalid),
    .dmem_arready(friscv_dmem_arready),
    .dmem_araddr(friscv_dmem_araddr),
    .dmem_arprot(friscv_dmem_arprot),
    .dmem_arid(friscv_dmem_arid),
    .dmem_rvalid(friscv_dmem_rvalid),
    .dmem_rready(friscv_dmem_rready),
    .dmem_rid(friscv_dmem_rid),
    .dmem_rresp(friscv_dmem_rresp),
    .dmem_rdata(friscv_dmem_rdata)
);

// ==============================================================================
// Width Adapter: Instruction Bus (128→32)
// ==============================================================================
axi_width_adapter_128to32 #(
    .MASTER_DATA_W(128),
    .SLAVE_DATA_W(32),
    .ADDR_W(32),
    .ID_W(8)
) u_instr_width_adapter (
    .aclk(ACLK),
    .aresetn(ARESETN),
    
    // Master side (from FRISCV 128-bit)
    .m_awvalid(1'b0),              // Instruction bus is read-only
    .m_awready(),
    .m_awaddr(32'h0),
    .m_awprot(3'h0),
    .m_awid(8'h0),
    .m_wvalid(1'b0),
    .m_wready(),
    .m_wdata(128'h0),
    .m_wstrb(16'h0),
    .m_bvalid(),
    .m_bready(1'b1),
    .m_bid(),
    .m_bresp(),
    
    .m_arvalid(friscv_imem_arvalid),
    .m_arready(friscv_imem_arready),
    .m_araddr(friscv_imem_araddr),
    .m_arprot(friscv_imem_arprot),
    .m_arid(friscv_imem_arid),
    .m_rvalid(friscv_imem_rvalid),
    .m_rready(friscv_imem_rready),
    .m_rid(friscv_imem_rid),
    .m_rresp(friscv_imem_rresp),
    .m_rdata(friscv_imem_rdata),
    
    // Slave side (to Interconnect 32-bit)
    .s_awvalid(),                  // Unused (read-only)
    .s_awready(1'b1),
    .s_awaddr(),
    .s_awprot(),
    .s_awid(),
    .s_wvalid(),
    .s_wready(1'b1),
    .s_wdata(),
    .s_wstrb(),
    .s_bvalid(1'b0),
    .s_bready(),
    .s_bid(8'h0),
    .s_bresp(2'b00),
    
    .s_arvalid(m0_axi_arvalid),
    .s_arready(m0_axi_arready),
    .s_araddr(m0_axi_araddr),
    .s_arprot(m0_axi_arprot),
    .s_arid(),                     // Not used by interconnect
    .s_rvalid(m0_axi_rvalid),
    .s_rready(m0_axi_rready),
    .s_rid(8'h0),
    .s_rresp(m0_axi_rresp),
    .s_rdata(m0_axi_rdata)
);

// ==============================================================================
// Width Adapter: Data Bus (128→32)
// ==============================================================================
axi_width_adapter_128to32 #(
    .MASTER_DATA_W(128),
    .SLAVE_DATA_W(32),
    .ADDR_W(32),
    .ID_W(8)
) u_data_width_adapter (
    .aclk(ACLK),
    .aresetn(ARESETN),
    
    // Master side (from FRISCV 128-bit)
    .m_awvalid(friscv_dmem_awvalid),
    .m_awready(friscv_dmem_awready),
    .m_awaddr(friscv_dmem_awaddr),
    .m_awprot(friscv_dmem_awprot),
    .m_awid(friscv_dmem_awid),
    .m_wvalid(friscv_dmem_wvalid),
    .m_wready(friscv_dmem_wready),
    .m_wdata(friscv_dmem_wdata),
    .m_wstrb(friscv_dmem_wstrb),
    .m_bvalid(friscv_dmem_bvalid),
    .m_bready(friscv_dmem_bready),
    .m_bid(friscv_dmem_bid),
    .m_bresp(friscv_dmem_bresp),
    .m_arvalid(friscv_dmem_arvalid),
    .m_arready(friscv_dmem_arready),
    .m_araddr(friscv_dmem_araddr),
    .m_arprot(friscv_dmem_arprot),
    .m_arid(friscv_dmem_arid),
    .m_rvalid(friscv_dmem_rvalid),
    .m_rready(friscv_dmem_rready),
    .m_rid(friscv_dmem_rid),
    .m_rresp(friscv_dmem_rresp),
    .m_rdata(friscv_dmem_rdata),
    
    // Slave side (to Interconnect 32-bit)
    .s_awvalid(m1_axi_awvalid),
    .s_awready(m1_axi_awready),
    .s_awaddr(m1_axi_awaddr),
    .s_awprot(m1_axi_awprot),
    .s_awid(),
    .s_wvalid(m1_axi_wvalid),
    .s_wready(m1_axi_wready),
    .s_wdata(m1_axi_wdata),
    .s_wstrb(m1_axi_wstrb),
    .s_bvalid(m1_axi_bvalid),
    .s_bready(m1_axi_bready),
    .s_bid(8'h0),
    .s_bresp(m1_axi_bresp),
    .s_arvalid(m1_axi_arvalid),
    .s_arready(m1_axi_arready),
    .s_araddr(m1_axi_araddr),
    .s_arprot(m1_axi_arprot),
    .s_arid(),
    .s_rvalid(m1_axi_rvalid),
    .s_rready(m1_axi_rready),
    .s_rid(8'h0),
    .s_rresp(m1_axi_rresp),
    .s_rdata(m1_axi_rdata)
);

// ==============================================================================
// AXI Interconnect (2M × 4S)
// ==============================================================================
// ==============================================================================
// AXI Interconnect - Using AXI_Interconnect_Full (supports 4 slaves)
// ==============================================================================
// Port Mapping:
//   S00_AXI_* = Master 0 (Instruction - Read only)
//   S01_AXI_* = Master 1 (Data - Read/Write)
//   M00_AXI_* = Slave 0 (RAM)
//   M01_AXI_* = Slave 1 (GPIO)
//   M02_AXI_* = Slave 2 (UART)
//   M03_AXI_* = Slave 3 (SPI)
// ==============================================================================

AXI_Interconnect_Full #(
    .ARBITRATION_MODE(1)  // Round-Robin
) u_axi_interconnect (
    .ACLK(ACLK),
    .ARESETN(ARESETN),
    
    // Slave address ranges
    .slave0_addr1(32'h00000000),  // RAM base
    .slave0_addr2(32'h1FFFFFFF),  // RAM end
    .slave1_addr1(32'h40000000),  // GPIO base
    .slave1_addr2(32'h5FFFFFFF),  // GPIO end
    .slave2_addr1(32'h80000000),  // UART base
    .slave2_addr2(32'hBFFFFFFF),  // UART end
    .slave3_addr1(32'hC0000000),  // SPI base
    .slave3_addr2(32'hFFFFFFFF),  // SPI end
    
    // ========================================================================
    // S00: Master 0 (Instruction - Read only)
    // ========================================================================
    .S00_ACLK(ACLK),
    .S00_ARESETN(ARESETN),
    // Write channels (unused - instruction is read-only)
    .S00_AXI_awaddr(32'h0),
    .S00_AXI_awlen(8'h0),
    .S00_AXI_awsize(3'h0),
    .S00_AXI_awburst(2'h0),
    .S00_AXI_awlock(2'h0),
    .S00_AXI_awcache(4'h0),
    .S00_AXI_awprot(3'h0),
    .S00_AXI_awqos(4'h0),
    .S00_AXI_awvalid(1'b0),
    .S00_AXI_awready(),
    .S00_AXI_wdata(32'h0),
    .S00_AXI_wstrb(4'h0),
    .S00_AXI_wlast(1'b0),
    .S00_AXI_wvalid(1'b0),
    .S00_AXI_wready(),
    .S00_AXI_bresp(),
    .S00_AXI_bvalid(),
    .S00_AXI_bready(1'b1),
    // Read channels
    .S00_AXI_araddr(m0_axi_araddr),
    .S00_AXI_arlen(8'h00),
    .S00_AXI_arsize(3'b010),
    .S00_AXI_arburst(2'b01),
    .S00_AXI_arlock(2'h0),
    .S00_AXI_arcache(4'h0),
    .S00_AXI_arprot(m0_axi_arprot),
    .S00_AXI_arregion(4'h0),
    .S00_AXI_arqos(4'h0),
    .S00_AXI_arvalid(m0_axi_arvalid),
    .S00_AXI_arready(m0_axi_arready),
    .S00_AXI_rdata(m0_axi_rdata),
    .S00_AXI_rresp(m0_axi_rresp),
    .S00_AXI_rlast(m0_axi_rlast),
    .S00_AXI_rvalid(m0_axi_rvalid),
    .S00_AXI_rready(m0_axi_rready),
    
    // ========================================================================
    // S01: Master 1 (Data - Read/Write)
    // ========================================================================
    .S01_ACLK(ACLK),
    .S01_ARESETN(ARESETN),
    // Write channels
    .S01_AXI_awaddr(m1_axi_awaddr),
    .S01_AXI_awlen(8'h00),
    .S01_AXI_awsize(3'b010),
    .S01_AXI_awburst(2'b01),
    .S01_AXI_awlock(2'h0),
    .S01_AXI_awcache(4'h0),
    .S01_AXI_awprot(m1_axi_awprot),
    .S01_AXI_awqos(4'h0),
    .S01_AXI_awvalid(m1_axi_awvalid),
    .S01_AXI_awready(m1_axi_awready),
    .S01_AXI_wdata(m1_axi_wdata),
    .S01_AXI_wstrb(m1_axi_wstrb),
    .S01_AXI_wlast(1'b1),
    .S01_AXI_wvalid(m1_axi_wvalid),
    .S01_AXI_wready(m1_axi_wready),
    .S01_AXI_bresp(m1_axi_bresp),
    .S01_AXI_bvalid(m1_axi_bvalid),
    .S01_AXI_bready(m1_axi_bready),
    // Read channels
    .S01_AXI_araddr(m1_axi_araddr),
    .S01_AXI_arlen(8'h00),
    .S01_AXI_arsize(3'b010),
    .S01_AXI_arburst(2'b01),
    .S01_AXI_arlock(2'h0),
    .S01_AXI_arcache(4'h0),
    .S01_AXI_arprot(m1_axi_arprot),
    .S01_AXI_arregion(4'h0),
    .S01_AXI_arqos(4'h0),
    .S01_AXI_arvalid(m1_axi_arvalid),
    .S01_AXI_arready(m1_axi_arready),
    .S01_AXI_rdata(m1_axi_rdata),
    .S01_AXI_rresp(m1_axi_rresp),
    .S01_AXI_rlast(m1_axi_rlast),
    .S01_AXI_rvalid(m1_axi_rvalid),
    .S01_AXI_rready(m1_axi_rready),
    
    // ========================================================================
    // M00: Slave 0 (RAM)
    // ========================================================================
    .M00_ACLK(ACLK),
    .M00_ARESETN(ARESETN),
    .M00_AXI_awaddr_ID(),  // Unused
    .M00_AXI_awaddr(s0_axi_awaddr),
    .M00_AXI_awlen(8'h00),
    .M00_AXI_awsize(3'b010),
    .M00_AXI_awburst(2'b01),
    .M00_AXI_awlock(),
    .M00_AXI_awcache(),
    .M00_AXI_awprot(),
    .M00_AXI_awqos(),
    .M00_AXI_awvalid(s0_axi_awvalid),
    .M00_AXI_awready(s0_axi_awready),
    .M00_AXI_wdata(s0_axi_wdata),
    .M00_AXI_wstrb(s0_axi_wstrb),
    .M00_AXI_wlast(1'b1),
    .M00_AXI_wvalid(s0_axi_wvalid),
    .M00_AXI_wready(s0_axi_wready),
    .M00_AXI_BID(1'b0),  // AXI-Lite doesn't use BID
    .M00_AXI_bresp(s0_axi_bresp),
    .M00_AXI_bvalid(s0_axi_bvalid),
    .M00_AXI_bready(s0_axi_bready),
    .M00_AXI_araddr(s0_axi_araddr),
    .M00_AXI_arlen(8'h00),
    .M00_AXI_arsize(3'b010),
    .M00_AXI_arburst(2'b01),
    .M00_AXI_arlock(),
    .M00_AXI_arcache(),
    .M00_AXI_arprot(),
    .M00_AXI_arregion(),
    .M00_AXI_arqos(),
    .M00_AXI_arvalid(s0_axi_arvalid),
    .M00_AXI_arready(s0_axi_arready),
    .M00_AXI_rdata(s0_axi_rdata),
    .M00_AXI_rresp(s0_axi_rresp),
    .M00_AXI_rlast(1'b1),
    .M00_AXI_rvalid(s0_axi_rvalid),
    .M00_AXI_rready(s0_axi_rready),
    
    // ========================================================================
    // M01: Slave 1 (GPIO)
    // ========================================================================
    .M01_ACLK(ACLK),
    .M01_ARESETN(ARESETN),
    .M01_AXI_awaddr_ID(),  // Unused
    .M01_AXI_awaddr(s1_axi_awaddr),
    .M01_AXI_awlen(8'h00),
    .M01_AXI_awsize(3'b010),
    .M01_AXI_awburst(2'b01),
    .M01_AXI_awlock(),
    .M01_AXI_awcache(),
    .M01_AXI_awprot(),
    .M01_AXI_awqos(),
    .M01_AXI_awvalid(s1_axi_awvalid),
    .M01_AXI_awready(s1_axi_awready),
    .M01_AXI_wdata(s1_axi_wdata),
    .M01_AXI_wstrb(s1_axi_wstrb),
    .M01_AXI_wlast(1'b1),
    .M01_AXI_wvalid(s1_axi_wvalid),
    .M01_AXI_wready(s1_axi_wready),
    .M01_AXI_BID(1'b0),
    .M01_AXI_bresp(s1_axi_bresp),
    .M01_AXI_bvalid(s1_axi_bvalid),
    .M01_AXI_bready(s1_axi_bready),
    .M01_AXI_araddr(s1_axi_araddr),
    .M01_AXI_arlen(8'h00),
    .M01_AXI_arsize(3'b010),
    .M01_AXI_arburst(2'b01),
    .M01_AXI_arlock(),
    .M01_AXI_arcache(),
    .M01_AXI_arprot(),
    .M01_AXI_arregion(),
    .M01_AXI_arqos(),
    .M01_AXI_arvalid(s1_axi_arvalid),
    .M01_AXI_arready(s1_axi_arready),
    .M01_AXI_rdata(s1_axi_rdata),
    .M01_AXI_rresp(s1_axi_rresp),
    .M01_AXI_rlast(1'b1),
    .M01_AXI_rvalid(s1_axi_rvalid),
    .M01_AXI_rready(s1_axi_rready),
    
    // ========================================================================
    // M02: Slave 2 (UART)
    // ========================================================================
    .M02_ACLK(ACLK),
    .M02_ARESETN(ARESETN),
    .M02_AXI_awaddr_ID(),  // Unused
    .M02_AXI_awaddr(s2_axi_awaddr),
    .M02_AXI_awlen(8'h00),
    .M02_AXI_awsize(3'b010),
    .M02_AXI_awburst(2'b01),
    .M02_AXI_awlock(),
    .M02_AXI_awcache(),
    .M02_AXI_awprot(),
    .M02_AXI_awqos(),
    .M02_AXI_awvalid(s2_axi_awvalid),
    .M02_AXI_awready(s2_axi_awready),
    .M02_AXI_wdata(s2_axi_wdata),
    .M02_AXI_wstrb(s2_axi_wstrb),
    .M02_AXI_wlast(1'b1),
    .M02_AXI_wvalid(s2_axi_wvalid),
    .M02_AXI_wready(s2_axi_wready),
    .M02_AXI_BID(1'b0),
    .M02_AXI_bresp(s2_axi_bresp),
    .M02_AXI_bvalid(s2_axi_bvalid),
    .M02_AXI_bready(s2_axi_bready),
    .M02_AXI_araddr(s2_axi_araddr),
    .M02_AXI_arlen(8'h00),
    .M02_AXI_arsize(3'b010),
    .M02_AXI_arburst(2'b01),
    .M02_AXI_arlock(),
    .M02_AXI_arcache(),
    .M02_AXI_arprot(),
    .M02_AXI_arregion(),
    .M02_AXI_arqos(),
    .M02_AXI_arvalid(s2_axi_arvalid),
    .M02_AXI_arready(s2_axi_arready),
    .M02_AXI_rdata(s2_axi_rdata),
    .M02_AXI_rresp(s2_axi_rresp),
    .M02_AXI_rlast(1'b1),
    .M02_AXI_rvalid(s2_axi_rvalid),
    .M02_AXI_rready(s2_axi_rready),
    
    // ========================================================================
    // M03: Slave 3 (SPI)
    // ========================================================================
    .M03_ACLK(ACLK),
    .M03_ARESETN(ARESETN),
    .M03_AXI_awaddr_ID(),  // Unused
    .M03_AXI_awaddr(s3_axi_awaddr),
    .M03_AXI_awlen(8'h00),
    .M03_AXI_awsize(3'b010),
    .M03_AXI_awburst(2'b01),
    .M03_AXI_awlock(),
    .M03_AXI_awcache(),
    .M03_AXI_awprot(),
    .M03_AXI_awqos(),
    .M03_AXI_awvalid(s3_axi_awvalid),
    .M03_AXI_awready(s3_axi_awready),
    .M03_AXI_wdata(s3_axi_wdata),
    .M03_AXI_wstrb(s3_axi_wstrb),
    .M03_AXI_wlast(1'b1),
    .M03_AXI_wvalid(s3_axi_wvalid),
    .M03_AXI_wready(s3_axi_wready),
    .M03_AXI_BID(1'b0),
    .M03_AXI_bresp(s3_axi_bresp),
    .M03_AXI_bvalid(s3_axi_bvalid),
    .M03_AXI_bready(s3_axi_bready),
    .M03_AXI_araddr(s3_axi_araddr),
    .M03_AXI_arlen(8'h00),
    .M03_AXI_arsize(3'b010),
    .M03_AXI_arburst(2'b01),
    .M03_AXI_arlock(),
    .M03_AXI_arcache(),
    .M03_AXI_arprot(),
    .M03_AXI_arregion(),
    .M03_AXI_arqos(),
    .M03_AXI_arvalid(s3_axi_arvalid),
    .M03_AXI_arready(s3_axi_arready),
    .M03_AXI_rdata(s3_axi_rdata),
    .M03_AXI_rresp(s3_axi_rresp),
    .M03_AXI_rlast(1'b1),
    .M03_AXI_rvalid(s3_axi_rvalid),
    .M03_AXI_rready(s3_axi_rready)
);

// ==============================================================================
// Peripherals (Unchanged from previous system)
// ==============================================================================

axi_lite_ram #(
    .ADDR_WIDTH(16),
    .DATA_WIDTH(32)
) u_ram (
    // ✅ FIXED: Correct port names
    .ACLK(ACLK),
    .ARESETN(ARESETN),
    .S_AXI_awaddr(s0_axi_awaddr[15:0]),
    .S_AXI_awprot(3'b000),
    .S_AXI_awvalid(s0_axi_awvalid),
    .S_AXI_awready(s0_axi_awready),
    .S_AXI_wdata(s0_axi_wdata),
    .S_AXI_wstrb(s0_axi_wstrb),
    .S_AXI_wvalid(s0_axi_wvalid),
    .S_AXI_wready(s0_axi_wready),
    .S_AXI_bresp(s0_axi_bresp),
    .S_AXI_bvalid(s0_axi_bvalid),
    .S_AXI_bready(s0_axi_bready),
    .S_AXI_araddr(s0_axi_araddr[15:0]),
    .S_AXI_arprot(3'b000),
    .S_AXI_arvalid(s0_axi_arvalid),
    .S_AXI_arready(s0_axi_arready),
    .S_AXI_rdata(s0_axi_rdata),
    .S_AXI_rresp(s0_axi_rresp),
    .S_AXI_rvalid(s0_axi_rvalid),
    .S_AXI_rlast(),              // Output
    .S_AXI_rready(s0_axi_rready)
);

axi_lite_gpio #(
    .ADDR_WIDTH(12),
    .DATA_WIDTH(32)
) u_gpio (
    // ✅ FIXED: Correct port names
    .ACLK(ACLK),
    .ARESETN(ARESETN),
    .S_AXI_awaddr(s1_axi_awaddr[11:0]),
    .S_AXI_awprot(3'b000),
    .S_AXI_awvalid(s1_axi_awvalid),
    .S_AXI_awready(s1_axi_awready),
    .S_AXI_wdata(s1_axi_wdata),
    .S_AXI_wstrb(s1_axi_wstrb),
    .S_AXI_wvalid(s1_axi_wvalid),
    .S_AXI_wready(s1_axi_wready),
    .S_AXI_bresp(s1_axi_bresp),
    .S_AXI_bvalid(s1_axi_bvalid),
    .S_AXI_bready(s1_axi_bready),
    .S_AXI_araddr(s1_axi_araddr[11:0]),
    .S_AXI_arprot(3'b000),
    .S_AXI_arvalid(s1_axi_arvalid),
    .S_AXI_arready(s1_axi_arready),
    .S_AXI_rdata(s1_axi_rdata),
    .S_AXI_rresp(s1_axi_rresp),
    .S_AXI_rvalid(s1_axi_rvalid),
    .S_AXI_rlast(),              // Output
    .S_AXI_rready(s1_axi_rready),
    .gpio_in(gpio_in),
    .gpio_out(gpio_out)
);

axi_lite_uart #(
    .ADDR_WIDTH(12),
    .DATA_WIDTH(32)
) u_uart (
    // ✅ FIXED: Correct port names
    .ACLK(ACLK),
    .ARESETN(ARESETN),
    .S_AXI_awaddr(s2_axi_awaddr[11:0]),
    .S_AXI_awprot(3'b000),
    .S_AXI_awvalid(s2_axi_awvalid),
    .S_AXI_awready(s2_axi_awready),
    .S_AXI_wdata(s2_axi_wdata),
    .S_AXI_wstrb(s2_axi_wstrb),
    .S_AXI_wvalid(s2_axi_wvalid),
    .S_AXI_wready(s2_axi_wready),
    .S_AXI_bresp(s2_axi_bresp),
    .S_AXI_bvalid(s2_axi_bvalid),
    .S_AXI_bready(s2_axi_bready),
    .S_AXI_araddr(s2_axi_araddr[11:0]),
    .S_AXI_arprot(3'b000),
    .S_AXI_arvalid(s2_axi_arvalid),
    .S_AXI_arready(s2_axi_arready),
    .S_AXI_rdata(s2_axi_rdata),
    .S_AXI_rresp(s2_axi_rresp),
    .S_AXI_rvalid(s2_axi_rvalid),
    .S_AXI_rlast(),              // Output, not connected
    .S_AXI_rready(s2_axi_rready),
    .tx_valid(),                 // UART TX signals (not used in this system)
    .tx_byte()
);

axi_lite_spi #(
    .ADDR_WIDTH(12),
    .DATA_WIDTH(32)
) u_spi (
    // ✅ FIXED: Correct port names
    .ACLK(ACLK),
    .ARESETN(ARESETN),
    .S_AXI_awaddr(s3_axi_awaddr[11:0]),
    .S_AXI_awprot(3'b000),
    .S_AXI_awvalid(s3_axi_awvalid),
    .S_AXI_awready(s3_axi_awready),
    .S_AXI_wdata(s3_axi_wdata),
    .S_AXI_wstrb(s3_axi_wstrb),
    .S_AXI_wvalid(s3_axi_wvalid),
    .S_AXI_wready(s3_axi_wready),   // ✅ FIXED: was S3_AXI_wready
    .S_AXI_bresp(s3_axi_bresp),
    .S_AXI_bvalid(s3_axi_bvalid),
    .S_AXI_bready(s3_axi_bready),
    .S_AXI_araddr(s3_axi_araddr[11:0]),
    .S_AXI_arprot(3'b000),
    .S_AXI_arvalid(s3_axi_arvalid),
    .S_AXI_arready(s3_axi_arready),
    .S_AXI_rdata(s3_axi_rdata),
    .S_AXI_rresp(s3_axi_rresp),
    .S_AXI_rvalid(s3_axi_rvalid),
    .S_AXI_rlast(),              // Output, not connected
    .S_AXI_rready(s3_axi_rready),
    .spi_cs_n(spi_cs_n),
    .spi_sclk(spi_sclk),
    .spi_mosi(spi_mosi),
    .spi_miso(spi_miso)
);

endmodule

