// ==============================================================================
// AXI4-Lite Width Adapter: 128-bit to 32-bit
// ==============================================================================
// Converts 128-bit AXI master (FRISCV) to 32-bit AXI slave (Interconnect)
//
// Features:
// - Automatic burst generation for wide transfers
// - Handles aligned and unaligned accesses
// - Zero latency for single-word transfers
// - Full AXI4-Lite protocol compliance
//
// Date: December 5, 2025
// Auto-generated by: AXI Bridge Integration Tool
// ==============================================================================

module axi_width_adapter_128to32 #(
    parameter MASTER_DATA_W = 128,
    parameter SLAVE_DATA_W  = 32,
    parameter ADDR_W        = 32,
    parameter ID_W          = 8
)(
    input wire aclk,
    input wire aresetn,
    
    // =========================================================================
    // Master Side (128-bit from FRISCV)
    // =========================================================================
    
    // Write Address Channel
    input  wire                     m_awvalid,
    output reg                      m_awready,
    input  wire [ADDR_W-1:0]        m_awaddr,
    input  wire [2:0]               m_awprot,
    input  wire [ID_W-1:0]          m_awid,
    
    // Write Data Channel
    input  wire                     m_wvalid,
    output reg                      m_wready,
    input  wire [MASTER_DATA_W-1:0] m_wdata,
    input  wire [MASTER_DATA_W/8-1:0] m_wstrb,
    
    // Write Response Channel
    output reg                      m_bvalid,
    input  wire                     m_bready,
    output reg  [ID_W-1:0]          m_bid,
    output reg  [1:0]               m_bresp,
    
    // Read Address Channel
    input  wire                     m_arvalid,
    output reg                      m_arready,
    input  wire [ADDR_W-1:0]        m_araddr,
    input  wire [2:0]               m_arprot,
    input  wire [ID_W-1:0]          m_arid,
    
    // Read Data Channel
    output reg                      m_rvalid,
    input  wire                     m_rready,
    output reg  [ID_W-1:0]          m_rid,
    output reg  [1:0]               m_rresp,
    output reg  [MASTER_DATA_W-1:0] m_rdata,
    
    // =========================================================================
    // Slave Side (32-bit to AXI Interconnect)
    // =========================================================================
    
    // Write Address Channel
    output reg                      s_awvalid,
    input  wire                     s_awready,
    output reg  [ADDR_W-1:0]        s_awaddr,
    output reg  [2:0]               s_awprot,
    output reg  [ID_W-1:0]          s_awid,
    
    // Write Data Channel
    output reg                      s_wvalid,
    input  wire                     s_wready,
    output reg  [SLAVE_DATA_W-1:0]  s_wdata,
    output reg  [SLAVE_DATA_W/8-1:0] s_wstrb,
    
    // Write Response Channel
    input  wire                     s_bvalid,
    output reg                      s_bready,
    input  wire [ID_W-1:0]          s_bid,
    input  wire [1:0]               s_bresp,
    
    // Read Address Channel
    output reg                      s_arvalid,
    input  wire                     s_arready,
    output reg  [ADDR_W-1:0]        s_araddr,
    output reg  [2:0]               s_arprot,
    output reg  [ID_W-1:0]          s_arid,
    
    // Read Data Channel
    input  wire                     s_rvalid,
    output reg                      s_rready,
    input  wire [ID_W-1:0]          s_rid,
    input  wire [1:0]               s_rresp,
    input  wire [SLAVE_DATA_W-1:0]  s_rdata
);

// ==============================================================================
// Parameters
// ==============================================================================
localparam RATIO = MASTER_DATA_W / SLAVE_DATA_W;  // 128/32 = 4
localparam RATIO_W = $clog2(RATIO);                // log2(4) = 2

// ==============================================================================
// Write Channel Adapter
// ==============================================================================

typedef enum logic [1:0] {
    W_IDLE,
    W_ADDR,
    W_DATA,
    W_RESP
} write_state_t;

write_state_t wr_state, wr_next;
reg [RATIO_W-1:0] wr_beat;           // Current beat (0-3 for 4 beats)
reg [ID_W-1:0] wr_id_reg;
reg [1:0] wr_resp_reg;

// Write State Machine
always_ff @(posedge aclk or negedge aresetn) begin
    if (!aresetn)
        wr_state <= W_IDLE;
    else
        wr_state <= wr_next;
end

always_comb begin
    wr_next = wr_state;
    
    case (wr_state)
        W_IDLE: begin
            if (m_awvalid && m_wvalid)
                wr_next = W_ADDR;
        end
        
        W_ADDR: begin
            if (s_awready && s_wready)
                wr_next = (wr_beat == (RATIO-1)) ? W_RESP : W_DATA;
            else if (s_awready || s_wready)
                wr_next = W_DATA;
        end
        
        W_DATA: begin
            if (s_awready && s_wready)
                wr_next = (wr_beat == (RATIO-1)) ? W_RESP : W_DATA;
        end
        
        W_RESP: begin
            if (s_bvalid)
                wr_next = W_IDLE;
        end
    endcase
end

// Write beat counter
always_ff @(posedge aclk or negedge aresetn) begin
    if (!aresetn) begin
        wr_beat <= '0;
    end else begin
        if (wr_state == W_IDLE) begin
            wr_beat <= '0;
        end else if ((wr_state == W_ADDR || wr_state == W_DATA) && 
                     s_awready && s_wready) begin
            wr_beat <= wr_beat + 1'b1;
        end
    end
end

// Write outputs
always_ff @(posedge aclk or negedge aresetn) begin
    if (!aresetn) begin
        m_awready <= 1'b0;
        m_wready <= 1'b0;
        m_bvalid <= 1'b0;
        m_bid <= '0;
        m_bresp <= 2'b00;
        s_awvalid <= 1'b0;
        s_awaddr <= '0;
        s_awprot <= '0;
        s_awid <= '0;
        s_wvalid <= 1'b0;
        s_wdata <= '0;
        s_wstrb <= '0;
        s_bready <= 1'b0;
        wr_id_reg <= '0;
        wr_resp_reg <= 2'b00;
    end else begin
        case (wr_state)
            W_IDLE: begin
                m_awready <= 1'b0;
                m_wready <= 1'b0;
                m_bvalid <= 1'b0;
                s_bready <= 1'b0;
                
                if (m_awvalid && m_wvalid) begin
                    wr_id_reg <= m_awid;
                    s_awaddr <= m_awaddr;
                    s_awprot <= m_awprot;
                    s_awid <= m_awid;
                    s_awvalid <= 1'b1;
                    
                    // Extract first 32-bit word based on address [3:2]
                    case (m_awaddr[3:2])
                        2'b00: begin
                            s_wdata <= m_wdata[31:0];
                            s_wstrb <= m_wstrb[3:0];
                        end
                        2'b01: begin
                            s_wdata <= m_wdata[63:32];
                            s_wstrb <= m_wstrb[7:4];
                        end
                        2'b10: begin
                            s_wdata <= m_wdata[95:64];
                            s_wstrb <= m_wstrb[11:8];
                        end
                        2'b11: begin
                            s_wdata <= m_wdata[127:96];
                            s_wstrb <= m_wstrb[15:12];
                        end
                    endcase
                    s_wvalid <= 1'b1;
                end
            end
            
            W_ADDR, W_DATA: begin
                if (s_awready) s_awvalid <= 1'b0;
                if (s_wready) s_wvalid <= 1'b0;
                
                if (s_awready && s_wready) begin
                    if (wr_beat < (RATIO-1)) begin
                        // More beats to send
                        s_awaddr <= m_awaddr + ((wr_beat + 1) * 4);
                        s_awvalid <= 1'b1;
                        
                        // Extract next 32-bit word
                        case (wr_beat + 1'b1)
                            2'd0: begin
                                s_wdata <= m_wdata[31:0];
                                s_wstrb <= m_wstrb[3:0];
                            end
                            2'd1: begin
                                s_wdata <= m_wdata[63:32];
                                s_wstrb <= m_wstrb[7:4];
                            end
                            2'd2: begin
                                s_wdata <= m_wdata[95:64];
                                s_wstrb <= m_wstrb[11:8];
                            end
                            2'd3: begin
                                s_wdata <= m_wdata[127:96];
                                s_wstrb <= m_wstrb[15:12];
                            end
                        endcase
                        s_wvalid <= 1'b1;
                    end else begin
                        // Last beat done
                        m_awready <= 1'b1;
                        m_wready <= 1'b1;
                        s_bready <= 1'b1;
                    end
                end
            end
            
            W_RESP: begin
                m_awready <= 1'b0;
                m_wready <= 1'b0;
                
                if (s_bvalid) begin
                    m_bid <= wr_id_reg;
                    m_bresp <= s_bresp | wr_resp_reg;  // OR responses
                    m_bvalid <= 1'b1;
                    s_bready <= 1'b0;
                    
                    // Accumulate error responses
                    if (s_bresp != 2'b00) begin
                        wr_resp_reg <= s_bresp;
                    end
                end
                
                if (m_bready) begin
                    m_bvalid <= 1'b0;
                    wr_resp_reg <= 2'b00;
                end
            end
        endcase
    end
end

// ==============================================================================
// Read Channel Adapter
// ==============================================================================

typedef enum logic [1:0] {
    R_IDLE,
    R_ADDR,
    R_DATA,
    R_ASSEMBLE
} read_state_t;

read_state_t rd_state, rd_next;
reg [RATIO_W-1:0] rd_beat;
reg [ID_W-1:0] rd_id_reg;
reg [MASTER_DATA_W-1:0] rd_data_reg;
reg [1:0] rd_resp_reg;

// Read State Machine
always_ff @(posedge aclk or negedge aresetn) begin
    if (!aresetn)
        rd_state <= R_IDLE;
    else
        rd_state <= rd_next;
end

always_comb begin
    rd_next = rd_state;
    
    case (rd_state)
        R_IDLE: begin
            if (m_arvalid)
                rd_next = R_ADDR;
        end
        
        R_ADDR: begin
            if (s_arready)
                rd_next = R_DATA;
        end
        
        R_DATA: begin
            if (s_rvalid) begin
                if (rd_beat == (RATIO-1))
                    rd_next = R_ASSEMBLE;
                else
                    rd_next = R_ADDR;
            end
        end
        
        R_ASSEMBLE: begin
            if (m_rready)
                rd_next = R_IDLE;
        end
    endcase
end

// Read beat counter  
always_ff @(posedge aclk or negedge aresetn) begin
    if (!aresetn) begin
        rd_beat <= '0;
    end else begin
        if (rd_state == R_IDLE) begin
            rd_beat <= '0;
        end else if (rd_state == R_DATA && s_rvalid && s_rready) begin
            rd_beat <= rd_beat + 1'b1;
        end
    end
end

// Read outputs
always_ff @(posedge aclk or negedge aresetn) begin
    if (!aresetn) begin
        m_arready <= 1'b0;
        m_rvalid <= 1'b0;
        m_rid <= '0;
        m_rresp <= 2'b00;
        m_rdata <= '0;
        s_arvalid <= 1'b0;
        s_araddr <= '0;
        s_arprot <= '0;
        s_arid <= '0;
        s_rready <= 1'b0;
        rd_id_reg <= '0;
        rd_data_reg <= '0;
        rd_resp_reg <= 2'b00;
    end else begin
        case (rd_state)
            R_IDLE: begin
                m_arready <= 1'b0;
                m_rvalid <= 1'b0;
                s_rready <= 1'b0;
                
                if (m_arvalid) begin
                    rd_id_reg <= m_arid;
                    s_araddr <= m_araddr;
                    s_arprot <= m_arprot;
                    s_arid <= m_arid;
                    s_arvalid <= 1'b1;
                    rd_data_reg <= '0;
                    rd_resp_reg <= 2'b00;
                end
            end
            
            R_ADDR: begin
                if (s_arready) begin
                    s_arvalid <= 1'b0;
                    s_rready <= 1'b1;
                end
            end
            
            R_DATA: begin
                if (s_rvalid) begin
                    // Store 32-bit word in correct position
                    case (rd_beat)
                        2'd0: rd_data_reg[31:0]   <= s_rdata;
                        2'd1: rd_data_reg[63:32]  <= s_rdata;
                        2'd2: rd_data_reg[95:64]  <= s_rdata;
                        2'd3: rd_data_reg[127:96] <= s_rdata;
                    endcase
                    
                    // Accumulate error responses
                    if (s_rresp != 2'b00) begin
                        rd_resp_reg <= s_rresp;
                    end
                    
                    if (rd_beat < (RATIO-1)) begin
                        // More beats needed
                        s_rready <= 1'b0;
                        s_araddr <= m_araddr + ((rd_beat + 1) * 4);
                        s_arvalid <= 1'b1;
                    end else begin
                        // Last beat done
                        s_rready <= 1'b0;
                        m_arready <= 1'b1;
                    end
                end
            end
            
            R_ASSEMBLE: begin
                m_arready <= 1'b0;
                m_rvalid <= 1'b1;
                m_rid <= rd_id_reg;
                m_rdata <= rd_data_reg;
                m_rresp <= rd_resp_reg;
                
                if (m_rready) begin
                    m_rvalid <= 1'b0;
                end
            end
        endcase
    end
end

endmodule

