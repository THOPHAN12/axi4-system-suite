library verilog;
use verilog.vl_types.all;
entity Read_Addr_Channel_Dec is
    generic(
        Num_OF_Masters  : integer := 2;
        Masters_ID_Size : vl_notype;
        Address_width   : integer := 32;
        AXI4_AR_len     : integer := 8;
        Num_Of_Slaves   : integer := 4;
        Base_Addr_Width : vl_notype
    );
    port(
        Master_AXI_araddr_ID: in     vl_logic_vector;
        Master_AXI_araddr: in     vl_logic_vector;
        Master_AXI_arlen: in     vl_logic_vector;
        Master_AXI_arsize: in     vl_logic_vector(2 downto 0);
        Master_AXI_arburst: in     vl_logic_vector(1 downto 0);
        Master_AXI_arlock: in     vl_logic_vector(1 downto 0);
        Master_AXI_arcache: in     vl_logic_vector(3 downto 0);
        Master_AXI_arprot: in     vl_logic_vector(2 downto 0);
        Master_AXI_arqos: in     vl_logic_vector(3 downto 0);
        Master_AXI_arregion: in     vl_logic_vector(3 downto 0);
        Master_AXI_arvalid: in     vl_logic;
        M00_AXI_araddr_ID: out    vl_logic_vector;
        M00_AXI_araddr  : out    vl_logic_vector;
        M00_AXI_arlen   : out    vl_logic_vector;
        M00_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M00_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M00_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M00_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M00_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M00_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M00_AXI_arvalid : out    vl_logic;
        M00_AXI_arready : in     vl_logic;
        M01_AXI_araddr_ID: out    vl_logic_vector;
        M01_AXI_araddr  : out    vl_logic_vector;
        M01_AXI_arlen   : out    vl_logic_vector;
        M01_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M01_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M01_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M01_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M01_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M01_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M01_AXI_arvalid : out    vl_logic;
        M01_AXI_arready : in     vl_logic;
        M02_AXI_araddr_ID: out    vl_logic_vector;
        M02_AXI_araddr  : out    vl_logic_vector;
        M02_AXI_arlen   : out    vl_logic_vector;
        M02_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M02_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M02_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M02_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M02_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M02_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M02_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M02_AXI_arvalid : out    vl_logic;
        M02_AXI_arready : in     vl_logic;
        M03_AXI_araddr_ID: out    vl_logic_vector;
        M03_AXI_araddr  : out    vl_logic_vector;
        M03_AXI_arlen   : out    vl_logic_vector;
        M03_AXI_arsize  : out    vl_logic_vector(2 downto 0);
        M03_AXI_arburst : out    vl_logic_vector(1 downto 0);
        M03_AXI_arlock  : out    vl_logic_vector(1 downto 0);
        M03_AXI_arcache : out    vl_logic_vector(3 downto 0);
        M03_AXI_arprot  : out    vl_logic_vector(2 downto 0);
        M03_AXI_arregion: out    vl_logic_vector(3 downto 0);
        M03_AXI_arqos   : out    vl_logic_vector(3 downto 0);
        M03_AXI_arvalid : out    vl_logic;
        M03_AXI_arready : in     vl_logic;
        Sel_Slave_Ready : out    vl_logic;
        Q_Enables       : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of Num_OF_Masters : constant is 1;
    attribute mti_svvh_generic_type of Masters_ID_Size : constant is 3;
    attribute mti_svvh_generic_type of Address_width : constant is 1;
    attribute mti_svvh_generic_type of AXI4_AR_len : constant is 1;
    attribute mti_svvh_generic_type of Num_Of_Slaves : constant is 1;
    attribute mti_svvh_generic_type of Base_Addr_Width : constant is 3;
end Read_Addr_Channel_Dec;
