//==============================================================================
// tb_arbitration_test.v
// Testbench for AXI Interconnect Arbitration Testing
//
// Tests 3 arbitration modes:
//   - Mode 0: FIXED_PRIORITY (Master 0 always wins)
//   - Mode 1: ROUND_ROBIN (Fair alternating - DEFAULT)
//   - Mode 2: QOS_BASED (Higher QoS value wins)
//
// Creates contention scenarios where both masters request simultaneously
//==============================================================================

`timescale 1ns/1ps

module tb_arbitration_test;

    //==========================================================================
    // Parameters
    //==========================================================================
    parameter ADDR_WIDTH = 32;
    parameter DATA_WIDTH = 32;
    parameter ID_WIDTH = 4;
    parameter RAM_WORDS = 2048;
    parameter CLK_PERIOD = 20;
    
    // Test configuration
    integer test_mode = 0;  // Will test modes 0, 1, 2
    
    //==========================================================================
    // Signals
    //==========================================================================
    reg ACLK;
    reg ARESETN;
    reg serv0_timer_irq;
    reg serv1_timer_irq;
    reg [31:0] gpio_in;
    reg spi_miso;
    
    wire [31:0] gpio_out;
    wire uart_tx_valid;
    wire [7:0] uart_tx_byte;
    wire spi_cs_n;
    wire spi_sclk;
    wire spi_mosi;
    
    //==========================================================================
    // Counters
    //==========================================================================
    integer m0_write_grants = 0;
    integer m1_write_grants = 0;
    integer m0_read_grants = 0;
    integer m1_read_grants = 0;
    
    //==========================================================================
    // DUT Instantiation - Will be recreated for each test mode
    //==========================================================================
    // Note: We'll need to use defparam or restart simulation for different modes
    // For now, using default mode (Round-Robin)
    
    dual_riscv_axi_system #(
        .ADDR_WIDTH  (ADDR_WIDTH),
        .DATA_WIDTH  (DATA_WIDTH),
        .ID_WIDTH    (ID_WIDTH),
        .RAM_WORDS   (RAM_WORDS),
        .RAM_INIT_HEX("")  // No program needed
    ) dut (
        .ACLK           (ACLK),
        .ARESETN        (ARESETN),
        .serv0_timer_irq(serv0_timer_irq),
        .serv1_timer_irq(serv1_timer_irq),
        .gpio_in        (gpio_in),
        .gpio_out       (gpio_out),
        .uart_tx_valid  (uart_tx_valid),
        .uart_tx_byte   (uart_tx_byte),
        .spi_cs_n       (spi_cs_n),
        .spi_sclk       (spi_sclk),
        .spi_mosi       (spi_mosi),
        .spi_miso       (spi_miso)
    );
    
    //==========================================================================
    // Clock Generation
    //==========================================================================
    initial begin
        ACLK = 0;
        forever #(CLK_PERIOD/2) ACLK = ~ACLK;
    end
    
    //==========================================================================
    // Banner
    //==========================================================================
    initial begin
        $display("\n//////////////////////////////////////////////////////////////////");
        $display("/  ARBITRATION TEST - AXI Interconnect                          /");
        $display("//////////////////////////////////////////////////////////////////\n");
        $display(" Test Purpose: Verify arbitration when both masters");
        $display("               request simultaneously (contention)\n");
        $display(" Arbitration Modes:");
        $display("   Mode 0: FIXED_PRIORITY - Master 0 always wins");
        $display("   Mode 1: ROUND_ROBIN - Fair alternating (DEFAULT)");
        $display("   Mode 2: QOS_BASED - Higher QoS value wins\n");
        $display("//////////////////////////////////////////////////////////////////\n");
    end
    
    //==========================================================================
    // Monitor Arbitration Grants
    //==========================================================================
    
    // Monitor Write Arbitration
    always @(posedge ACLK) begin
        if (ARESETN) begin
            // Check grant signals
            if (dut.u_axi_interconnect.u_full_interconnect.grant_m0_write) begin
                $display("[%0t] WRITE GRANT → Master 0", $time);
                m0_write_grants = m0_write_grants + 1;
            end
            
            if (dut.u_axi_interconnect.u_full_interconnect.grant_m1_write) begin
                $display("[%0t] WRITE GRANT → Master 1", $time);
                m1_write_grants = m1_write_grants + 1;
            end
        end
    end
    
    // Monitor Read Arbitration
    always @(posedge ACLK) begin
        if (ARESETN) begin
            if (dut.u_axi_interconnect.u_full_interconnect.grant_m0_read) begin
                $display("[%0t] READ GRANT TO Master 0", $time);
                m0_read_grants = m0_read_grants + 1;
            end
            
            if (dut.u_axi_interconnect.u_full_interconnect.grant_m1_read) begin
                $display("[%0t] READ GRANT TO Master 1", $time);
                m1_read_grants = m1_read_grants + 1;
            end
        end
    end
    
    // Monitor Arbiter State (Round-Robin) - Track turn changes
    reg [1:0] prev_wr_turn = 0;
    reg [1:0] prev_rd_turn = 0;
    
    always @(posedge ACLK) begin
        if (ARESETN) begin
            // Only for Round-Robin mode
            if (dut.u_axi_interconnect.ARBITRATION_MODE == 1) begin
                if (dut.u_axi_interconnect.u_full_interconnect.wr_turn !== prev_wr_turn) begin
                    $display("[%0t] WR_TURN changed TO %0d", $time, 
                            dut.u_axi_interconnect.u_full_interconnect.wr_turn);
                    prev_wr_turn = dut.u_axi_interconnect.u_full_interconnect.wr_turn;
                end
                if (dut.u_axi_interconnect.u_full_interconnect.rd_turn !== prev_rd_turn) begin
                    $display("[%0t] RD_TURN changed TO %0d", $time,
                            dut.u_axi_interconnect.u_full_interconnect.rd_turn);
                    prev_rd_turn = dut.u_axi_interconnect.u_full_interconnect.rd_turn;
                end
            end
        end
    end
    
    //==========================================================================
    // Test Scenario 1: WRITE Contention
    //==========================================================================
    task test_write_contention;
        input [255:0] mode_name;
        integer i;
        begin
            $display("\n//////////////////////////////////////////////////////////////////");
            $display("/  TEST: WRITE Contention - %s", mode_name);
            $display("//////////////////////////////////////////////////////////////////\n");
            
            $display("  Scenario: Both masters request WRITE simultaneously\n");
            
            // Reset counters
            m0_write_grants = 0;
            m1_write_grants = 0;
            
            // Wait a bit
            #100;
            
            $display("  Creating contention: Forcing both masters to request...\n");
            
            // Force both masters to request write simultaneously
            for (i = 0; i < 10; i = i + 1) begin
                // Master 0 Write Request
                force dut.serv0_axi_awvalid = 1;
                force dut.serv0_axi_awaddr = 32'h00000100 + (i * 4);
                force dut.serv0_axi_wvalid = 1;
                force dut.serv0_axi_wdata = 32'hAAAA0000 + i;
                force dut.serv0_axi_bready = 1;
                
                // Master 1 Write Request (SAME TIME!)
                force dut.serv1_axi_awvalid = 1;
                force dut.serv1_axi_awaddr = 32'h00000200 + (i * 4);
                force dut.serv1_axi_wvalid = 1;
                force dut.serv1_axi_wdata = 32'hBBBB0000 + i;
                force dut.serv1_axi_bready = 1;
                
                $display("  [Request %0d] Both masters requesting WRITE:", i+1);
                $display("    M0: Addr=0x%08h Data=0x%08h", 32'h00000100 + (i*4), 32'hAAAA0000 + i);
                $display("    M1: Addr=0x%08h Data=0x%08h", 32'h00000200 + (i*4), 32'hBBBB0000 + i);
                
                // Wait for transaction
                #(CLK_PERIOD * 5);
                
                // Release
                release dut.serv0_axi_awvalid;
                release dut.serv0_axi_wvalid;
                release dut.serv1_axi_awvalid;
                release dut.serv1_axi_wvalid;
                
                #(CLK_PERIOD * 2);
            end
            
            // Report results
            $display("\n  ━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━━");
            $display("  Results:");
            $display("    Master 0 Write Grants: %0d", m0_write_grants);
            $display("    Master 1 Write Grants: %0d", m1_write_grants);
            
            // Analyze results based on mode
            if (dut.u_axi_interconnect.ARBITRATION_MODE == 0) begin
                // Fixed Priority: M0 should win all
                $display("\n  Expected (Fixed Priority): M0 wins all");
                if (m0_write_grants > m1_write_grants) begin
                    $display(" CORRECT: M0 won %0d times (M1: %0d)", m0_write_grants, m1_write_grants);
                end else begin
                    $display(" Unexpected: M0=%0d M1=%0d", m0_write_grants, m1_write_grants);
                end
            end else if (dut.u_axi_interconnect.ARBITRATION_MODE == 1) begin
                // Round-Robin: Should alternate fairly
                $display("\n  Expected (Round-Robin): ~50/50 split");
                if (m0_write_grants >= 4 && m1_write_grants >= 4) begin
                    $display(" CORRECT: Fair split (M0=%0d, M1=%0d)", m0_write_grants, m1_write_grants);
                end else begin
                    $display(" Imbalanced: M0=%0d M1=%0d", m0_write_grants, m1_write_grants);
                end
            end else if (dut.u_axi_interconnect.ARBITRATION_MODE == 2) begin
                // QoS-based: Higher QoS wins
                $display("\n  Expected (QoS-based): Depends on QoS values");
                $display("  Result: M0=%0d M1=%0d", m0_write_grants, m1_write_grants);
            end
            
            $display("\n");
        end
    endtask
    
    //==========================================================================
    // Test Scenario 2: READ Contention
    //==========================================================================
    task test_read_contention;
        input [255:0] mode_name;
        integer i;
        begin
            $display("\n//////////////////////////////////////////////////////////////////");
            $display("/  TEST: READ Contention - %s", mode_name);
            $display("//////////////////////////////////////////////////////////////////\n");
            
            $display("  Scenario: Both masters request READ simultaneously\n");
            
            // Reset counters
            m0_read_grants = 0;
            m1_read_grants = 0;
            
            #100;
            
            $display("  Creating contention: Forcing both masters to request...\n");
            
            // Force both masters to request read simultaneously
            for (i = 0; i < 10; i = i + 1) begin
                // Master 0 Read Request
                force dut.serv0_axi_arvalid = 1;
                force dut.serv0_axi_araddr = 32'h00000300 + (i * 4);
                force dut.serv0_axi_rready = 1;
                
                // Master 1 Read Request (SAME TIME!)
                force dut.serv1_axi_arvalid = 1;
                force dut.serv1_axi_araddr = 32'h00000400 + (i * 4);
                force dut.serv1_axi_rready = 1;
                
                $display("  [Request %0d] Both masters requesting READ:", i+1);
                $display("    M0: Addr=0x%08h", 32'h00000300 + (i*4));
                $display("    M1: Addr=0x%08h", 32'h00000400 + (i*4));
                
                // Wait for transaction
                #(CLK_PERIOD * 5);
                
                // Release
                release dut.serv0_axi_arvalid;
                release dut.serv1_axi_arvalid;
                
                #(CLK_PERIOD * 2);
            end
            
            // Report results
            $display("\n////////////////////////////////////////////////////////////");
            $display("  Results:");
            $display("    Master 0 Read Grants: %0d", m0_read_grants);
            $display("    Master 1 Read Grants: %0d", m1_read_grants);
            
            // Analyze
            if (dut.u_axi_interconnect.ARBITRATION_MODE == 0) begin
                $display("\n  Expected (Fixed Priority): M0 wins all");
                if (m0_read_grants > m1_read_grants) begin
                    $display(" CORRECT: M0 won %0d times (M1: %0d)", m0_read_grants, m1_read_grants);
                end else begin
                    $display(" Unexpected: M0=%0d M1=%0d", m0_read_grants, m1_read_grants);
                end
            end else if (dut.u_axi_interconnect.ARBITRATION_MODE == 1) begin
                $display("\n  Expected (Round-Robin): ~50/50 split");
                if (m0_read_grants >= 4 && m1_read_grants >= 4) begin
                    $display(" CORRECT: Fair split (M0=%0d, M1=%0d)", m0_read_grants, m1_read_grants);
                end else begin
                    $display(" Imbalanced: M0=%0d M1=%0d", m0_read_grants, m1_read_grants);
                end
            end else if (dut.u_axi_interconnect.ARBITRATION_MODE == 2) begin
                $display("\n  Expected (QoS-based): Depends on QoS values");
                $display("  Result: M0=%0d M1=%0d", m0_read_grants, m1_read_grants);
            end
            
            $display("\n");
        end
    endtask
    
    //==========================================================================
    // Main Test Sequence
    //==========================================================================
    initial begin
        // Initialize
        serv0_timer_irq = 0;
        serv1_timer_irq = 0;
        gpio_in = 32'h0;
        spi_miso = 0;
        ARESETN = 0;
        
        // Reset
        #(CLK_PERIOD * 5);
        ARESETN = 1;
        #(CLK_PERIOD * 2);
        
        $display("[%0t] ✓ Reset complete\n", $time);
        $display("  Current Arbitration Mode: %0d", dut.u_axi_interconnect.ARBITRATION_MODE);
        
        case (dut.u_axi_interconnect.ARBITRATION_MODE)
            0: $display("  Mode Name: FIXED_PRIORITY");
            1: $display("  Mode Name: ROUND_ROBIN (DEFAULT)");
            2: $display("  Mode Name: QOS_BASED");
            default: $display("  Mode Name: UNKNOWN");
        endcase
        
        $display("\n");
        
        //======================================================================
        // Run Contention Tests
        //======================================================================
        
        test_write_contention("Current Mode");
        test_read_contention("Current Mode");
        
        //======================================================================
        // Final Summary
        //======================================================================
        $display("\n//////////////////////////////////////////////////////////////////");
        $display("/                    ARBITRATION TEST SUMMARY                    /");
        $display("//////////////////////////////////////////////////////////////////\n");
        
        $display(" Arbitration Mode: %0d", dut.u_axi_interconnect.ARBITRATION_MODE);
        case (dut.u_axi_interconnect.ARBITRATION_MODE)
            0: $display(" Mode: FIXED_PRIORITY");
            1: $display(" Mode: ROUND_ROBIN");
            2: $display(" Mode: QOS_BASED");
        endcase
        
        $display("\n Total Grants:");
        $display("  ////////////////////////////////////////////////////////////////////");
        $display("  Write Channel:");
        $display("    Master 0: %0d grants", m0_write_grants);
        $display("    Master 1: %0d grants", m1_write_grants);
        $display("    Total:    %0d", m0_write_grants + m1_write_grants);
        
        $display("\n  Read Channel:");
        $display("    Master 0: %0d grants", m0_read_grants);
        $display("    Master 1: %0d grants", m1_read_grants);
        $display("    Total:    %0d", m0_read_grants + m1_read_grants);
        
        $display("\n  Grand Total: %0d grants", 
                m0_write_grants + m1_write_grants + m0_read_grants + m1_read_grants);
        
        // Verify arbitration behavior
        $display("\n Arbitration Behavior Analysis:");
        $display("  ////////////////////////////////////////////////////////////////////");
        
        if (dut.u_axi_interconnect.ARBITRATION_MODE == 1) begin
            // Round-Robin expectations - calculate differences
            $display("  Write difference: %0d (Should be is less than or equal to 2 for fair RR)", 
                    (m0_write_grants > m1_write_grants) ? 
                    (m0_write_grants - m1_write_grants) : 
                    (m1_write_grants - m0_write_grants));
            $display("  Read difference:  %0d (Should be is less than or equal to 2 for fair RR 2 for fair RR)", 
                    (m0_read_grants > m1_read_grants) ? 
                    (m0_read_grants - m1_read_grants) : 
                    (m1_read_grants - m0_read_grants));
            
            // Check fairness
            if ((m0_write_grants >= 4) && (m1_write_grants >= 4) &&
                (m0_read_grants >= 4) && (m1_read_grants >= 4)) begin
                $display("\n ROUND_ROBIN: Working correctly!");
                $display("  Fair arbitration confirmed");
            end else begin
                $display("\n Round-Robin may have issues");
            end
        end
        
        $display("\n//////////////////////////////////////////////////////////////////");
        $display("/                    TEST COMPLETE                               /");
        $display("//////////////////////////////////////////////////////////////////\n");
        
        $display(" Arbitration logic verified");
        $display(" Contention scenarios tested");
        $display(" Both Write and Read channels tested\n");
        
        $finish;
    end
    
    //==========================================================================
    // Timeout
    //==========================================================================
    initial begin
        #500000;  // 500us timeout
        $display("\n Test complete (timeout)\n");
        $finish;
    end

endmodule

